module top_module(
    input clk,
    input [7:0] in,
    input reset,    // Synchronous reset
    output done); //
    
	parameter A = 0, B = 1, C = 2, D = 3;
    reg [1:0] pstate, nstate;
    // State transition logic (combinational)
    always @(*)
        begin
            case(pstate)
                A:nstate=in[3]?B:A;
                B:nstate = C;
                C:nstate = D;
                D:nstate = in[3]?B:A;
            endcase
        end
    // State flip-flops (sequential)
    always @(posedge clk)
        begin
            if(reset)
                pstate<=A;
            else
                pstate<=nstate;
        end
 
    // Output logic
    assign done = (pstate == D);

endmodule
