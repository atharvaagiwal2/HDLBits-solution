module top_module (
    input in,
    output out);
    always @(*)
        begin
            out = in;
        end
endmodule
