module top_module( input in, output out );
assign out = in; 
  //wire is directional, this means information flows in only one direction, from (usually one) source to the sinks
endmodule
